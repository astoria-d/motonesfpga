
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_arith.all;
use std.textio.all;

entity testbench_chr_rom is
end testbench_chr_rom;

architecture stimulus of testbench_chr_rom is 

begin
end stimulus ;

