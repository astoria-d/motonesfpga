
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_arith.all;
use std.textio.all;

entity testbench_motones_sim is
end testbench_motones_sim;

architecture stimulus of testbench_motones_sim is 
    constant cpu_clk : time := 589 ns;
    constant dsize : integer := 8;

begin
end stimulus ;

