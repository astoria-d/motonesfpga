library ieee;
use ieee.std_logic_1164.all;

entity ppu is 
    port (  clk         : in std_logic;
            ce_n        : in std_logic;
            rst_n       : in std_logic;
            r_nw        : in std_logic;
            cpu_addr    : in std_logic_vector (2 downto 0);
            cpu_d       : inout std_logic_vector (7 downto 0);
            vblank_n    : out std_logic;
            rd_n        : out std_logic;
            wr_n        : out std_logic;
            ale         : out std_logic;
            vram_ad     : inout std_logic_vector (7 downto 0);
            vram_a      : out std_logic_vector (13 downto 8);
            vga_clk     : in std_logic;
            h_sync_n    : out std_logic;
            v_sync_n    : out std_logic;
            r           : out std_logic_vector(3 downto 0);
            g           : out std_logic_vector(3 downto 0);
            b           : out std_logic_vector(3 downto 0)
    );
end ppu;

architecture rtl of ppu is

component ppu_render
    port (  clk         : in std_logic;
            rst_n       : in std_logic;
            vblank_n    : out std_logic;
            rd_n        : out std_logic;
            wr_n        : out std_logic;
            ale         : out std_logic;
            vram_ad     : inout std_logic_vector (7 downto 0);
            vram_a      : out std_logic_vector (13 downto 8);
            pos_x       : out std_logic_vector (8 downto 0);
            pos_y       : out std_logic_vector (8 downto 0);
            r           : out std_logic_vector (3 downto 0);
            g           : out std_logic_vector (3 downto 0);
            b           : out std_logic_vector (3 downto 0);
            ppu_ctrl        : in std_logic_vector (7 downto 0);
            ppu_mask        : in std_logic_vector (7 downto 0);
            ppu_status      : out std_logic_vector (7 downto 0);
            ppu_scroll_x    : in std_logic_vector (7 downto 0);
            ppu_scroll_y    : in std_logic_vector (7 downto 0);
            r_nw            : in std_logic;
            oam_bus_ce_n    : in std_logic;
            oam_addr        : in std_logic_vector (7 downto 0);
            oam_data        : inout std_logic_vector (7 downto 0);
            plt_bus_ce_n    : in std_logic;
            plt_addr        : in std_logic_vector (4 downto 0);
            plt_data        : inout std_logic_vector (5 downto 0)
    );
end component;

component vga_ctl
    port (  ppu_clk     : in std_logic;
            vga_clk     : in std_logic;
            rst_n       : in std_logic;
            pos_x       : in std_logic_vector (8 downto 0);
            pos_y       : in std_logic_vector (8 downto 0);
            nes_r       : in std_logic_vector (3 downto 0);
            nes_g       : in std_logic_vector (3 downto 0);
            nes_b       : in std_logic_vector (3 downto 0);
            h_sync_n    : out std_logic;
            v_sync_n    : out std_logic;
            r           : out std_logic_vector(3 downto 0);
            g           : out std_logic_vector(3 downto 0);
            b           : out std_logic_vector(3 downto 0)
    );
end component;

component d_flip_flop
    generic (
            dsize : integer := 8
            );
    port (
            clk     : in std_logic;
            res_n   : in std_logic;
            set_n   : in std_logic;
            we_n    : in std_logic;
            d       : in std_logic_vector (dsize - 1 downto 0);
            q       : out std_logic_vector (dsize - 1 downto 0)
        );
end component;

component counter_register
    generic (
        dsize       : integer := 8
    );
    port (  clk         : in std_logic;
            rst_n       : in std_logic;
            set_n       : in std_logic;
            ce_n        : in std_logic;
            d           : in std_logic_vector(dsize - 1 downto 0);
            q           : out std_logic_vector(dsize - 1 downto 0)
    );
end component;

signal pos_x       : std_logic_vector (8 downto 0);
signal pos_y       : std_logic_vector (8 downto 0);
signal nes_r       : std_logic_vector (3 downto 0);
signal nes_g       : std_logic_vector (3 downto 0);
signal nes_b       : std_logic_vector (3 downto 0);

constant dsize     : integer := 8;

constant PPUCTRL   : std_logic_vector(2 downto 0) := "000";
constant PPUMASK   : std_logic_vector(2 downto 0) := "001";
constant PPUSTATUS : std_logic_vector(2 downto 0) := "010";
constant OAMADDR   : std_logic_vector(2 downto 0) := "011";
constant OAMDATA   : std_logic_vector(2 downto 0) := "100";
constant PPUSCROLL : std_logic_vector(2 downto 0) := "101";
constant PPUADDR   : std_logic_vector(2 downto 0) := "110";
constant PPUDATA   : std_logic_vector(2 downto 0) := "111";

signal clk_n            : std_logic;

signal ppu_ctrl_we_n    : std_logic;
signal ppu_mask_we_n    : std_logic;
signal ppu_status_we_n  : std_logic;
signal oam_bus_ce_n     : std_logic;
signal oam_addr_we_n    : std_logic;
signal oam_data_we_n    : std_logic;
signal ppu_scroll_x_we_n    : std_logic;
signal ppu_scroll_y_we_n    : std_logic;
signal ppu_scroll_cnt_ce_n  : std_logic;
signal ppu_addr_we_n        : std_logic;
signal ppu_addr_cnt_ce_n    : std_logic;
signal ppu_data_we_n    : std_logic;

signal ppu_ctrl         : std_logic_vector (dsize - 1 downto 0);
signal ppu_mask         : std_logic_vector (dsize - 1 downto 0);
signal ppu_status       : std_logic_vector (dsize - 1 downto 0);
signal oam_addr         : std_logic_vector (dsize - 1 downto 0);
signal oam_data         : std_logic_vector (dsize - 1 downto 0);
signal ppu_scroll_x     : std_logic_vector (dsize - 1 downto 0);
signal ppu_scroll_y     : std_logic_vector (dsize - 1 downto 0);
signal ppu_scroll_cnt   : std_logic_vector (0 downto 0);
signal ppu_addr         : std_logic_vector (13 downto 0);
signal ppu_addr_in      : std_logic_vector (13 downto 0);
signal ppu_addr_cnt     : std_logic_vector (0 downto 0);
signal ppu_data         : std_logic_vector (dsize - 1 downto 0);

signal plt_bus_ce_n     : std_logic;
signal plt_addr         : std_logic_vector (4 downto 0);
signal plt_data         : std_logic_vector (5 downto 0);

begin

    render_inst : ppu_render port map (clk, rst_n, vblank_n, 
            rd_n, wr_n, ale, vram_ad, vram_a,
            pos_x, pos_y, nes_r, nes_g, nes_b,
            ppu_ctrl, ppu_mask, ppu_status, ppu_scroll_x, ppu_scroll_y,
            r_nw, oam_bus_ce_n, oam_addr, oam_data,
            plt_bus_ce_n, plt_addr, plt_data);

--    render_ad_buf : tri_state_buffer generic map (dsize)
--            port map ('0', render_vram_ad, vram_ad);
--    render_d_buf : tri_state_buffer generic map (6)
--            port map ('0', render_vram_a, vram_a);

    vga_inst : vga_ctl port map (clk, vga_clk, rst_n, 
            pos_x, pos_y, nes_r, nes_g, nes_b,
            h_sync_n, v_sync_n, r, g, b);

    --PPU registers.
    clk_n <= not clk;
    ppu_ctrl_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', ppu_ctrl_we_n, cpu_d, ppu_ctrl);

    ppu_mask_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', ppu_mask_we_n, cpu_d, ppu_mask);

    ppu_status_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', ppu_status_we_n, cpu_d, ppu_status);

    oma_addr_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', oam_addr_we_n, cpu_d, oam_addr);
    oma_data_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', oam_data_we_n, cpu_d, oam_data);

    ppu_scroll_x_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', ppu_scroll_x_we_n, cpu_d, ppu_scroll_x);
    ppu_scroll_y_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', ppu_scroll_y_we_n, cpu_d, ppu_scroll_y);
    ppu_scroll_cnt_inst : counter_register generic map (1)
            port map (clk_n, rst_n, '1', ppu_scroll_cnt_ce_n, (others => '0'), ppu_scroll_cnt);

    ppu_addr_inst : d_flip_flop generic map(14)
            port map (clk_n, rst_n, '1', ppu_addr_we_n, ppu_addr_in, ppu_addr);
    ppu_addr_cnt_inst : counter_register generic map (1)
            port map (clk_n, rst_n, '1', ppu_addr_cnt_ce_n, (others => '0'), ppu_addr_cnt);
    ppu_data_inst : d_flip_flop generic map(dsize)
            port map (clk_n, rst_n, '1', ppu_data_we_n, cpu_d, ppu_data);


    clock_p : process (clk)
    begin

        if (clk'event and clk = '1') then
            if (ce_n = '0') then
                --register set.
                if(cpu_addr = PPUCTRL) then
                    ppu_ctrl_we_n <= '0';
                else
                    ppu_ctrl_we_n <= '1';
                end if;

                if(cpu_addr = PPUMASK) then
                    ppu_mask_we_n <= '0';
                else
                    ppu_mask_we_n <= '1';
                end if;

                if(cpu_addr = PPUSTATUS) then
                    ppu_status_we_n <= '0';
                else
                    ppu_status_we_n <= '1';
                end if;

                if(cpu_addr = OAMADDR) then
                    oam_addr_we_n <= '0';
                else
                    oam_addr_we_n <= '1';
                end if;

                if(cpu_addr = OAMDATA) then
                    oam_data_we_n <= '0';
                else
                    oam_data_we_n <= '1';
                end if;

                if(cpu_addr = PPUSCROLL) then
                    ppu_scroll_cnt_ce_n <= '0';
                    if (ppu_scroll_cnt(0) = '0') then
                        ppu_scroll_x_we_n <= '0';
                        ppu_scroll_y_we_n <= '1';
                    else
                        ppu_scroll_y_we_n <= '0';
                        ppu_scroll_x_we_n <= '1';
                    end if;
                else
                    ppu_scroll_x_we_n <= '1';
                    ppu_scroll_y_we_n <= '1';
                    ppu_scroll_cnt_ce_n <= '1';
                end if;

                if(cpu_addr = PPUADDR) then
                    ppu_addr_cnt_ce_n <= '0';
                    ppu_addr_we_n <= '0';
                    if (ppu_addr_cnt(0) = '0') then
                        ppu_addr_in <= cpu_d(5 downto 0) & ppu_addr(7 downto 0);
                        ale <= '1';
                    else
                        ppu_addr_in <= ppu_addr(13 downto 8) & cpu_d;
                        vram_ad <= ppu_addr(7 downto 0);
                        vram_a <= ppu_addr(13 downto 8);
                        ale <= '0';
                    end if;
                else
                    ppu_addr_cnt_ce_n <= '1';
                    ppu_addr_we_n <= '1';
                    ale <= '1';
                end if;

                if(cpu_addr = PPUDATA) then
                    ppu_data_we_n <= '0';
                    rd_n <= not r_nw;
                    wr_n <= r_nw;
                else
                    ppu_data_we_n <= '1';
                    rd_n <= '1';
                    wr_n <= '1';
                end if;

            else
                ppu_ctrl_we_n    <= '1';
                ppu_mask_we_n    <= '1';
                ppu_status_we_n  <= '1';
                oam_bus_ce_n     <= '1';
                oam_addr_we_n    <= '1';
                oam_data_we_n    <= '1';
                ppu_scroll_x_we_n    <= '1';
                ppu_scroll_y_we_n    <= '1';
                ppu_scroll_cnt_ce_n  <= '1';
                ppu_addr_we_n        <= '1';
                ppu_addr_cnt_ce_n    <= '1';
                ppu_data_we_n    <= '1';

                ale <= 'Z';
                rd_n <= 'Z';
                wr_n <= 'Z';
                vram_ad <= (others => 'Z');
                vram_a <= (others => 'Z');
            end if; --if (ce_n = '0') then
        else

        end if;--if (clk'event and clk = '1') then

    end process;

----test init value set.
--    p_palette_init : process
--    variable i : integer := 0;
--use ieee.std_logic_arith.all;
--constant ppu_clk_time : time := 186 ns;
--    begin
--        wait for 7 us;
--
--        --fill palette teble.
--        plt_bus_ce_n <= '0';
--        plt_r_nw <= '0';
--        for i in 0 to 32 loop
--            plt_addr <= conv_std_logic_vector(i, 5);
--            plt_data <= conv_std_logic_vector((i - 1) * 4 + 17, 6);
--            wait for ppu_clk_time;
--        end loop;
--        plt_bus_ce_n <= '1';
--
--        ---TODO: for the time being...
--        plt_bus_ce_n <= 'Z';
--        plt_r_nw <= 'Z';
--        plt_addr <= (others => 'Z');
--        plt_data <= (others => 'Z');
--
--        wait;
--    end process;

end rtl;

